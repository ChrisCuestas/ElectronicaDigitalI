`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// University: Universidad Nacional de Colombia
// Students: Christian Camilo Cuestas  Ibanez y Eliana Ortiz García 
// 
// Create Date:    08/05/2018 
// Module Name:     LCDmult
// Project Name:  Proyecto Digital I: Reloj de Ajedrez
// Target Devices: Nexys 4
// Description:
//
//////////////////////////////////////////////////////////////////////////////////
module LCDmult(
	input clk,
	input wire [5:0] min1,
	input wire [5:0] seg1,
	input wire [5:0] min2,
	input wire [5:0] seg2,
	output wire	[5:0]	lcd
    );



endmodule
