`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// University: Universidad Nacional de Colombia
// Students: Christian Camilo Cuestas  Ibanez y Eliana Ortiz García 
// 
// Create Date:    08/05/2018 
// Module Name:    LCDcontrol 
// Project Name:  Proyecto Digital I: Reloj de Ajedrez
// Target Devices: Nexys 4
// Description:
//
//////////////////////////////////////////////////////////////////////////////////
module LCDcontrol(
	input	wire				clk,
	input	wire				setTime,
	input	wire	[5:0]	timeIn,
	input	wire	[23:0]	countedTime,
	output wire	[5:0]			lcd
    );


endmodule
